`include "include/timescale.v"

module or1200_vlx_dp(/*AUTOARG*/

   );

 //high when a byte should be stored

endmodule // or1200_vlx_dp
// Local Variables:
// verilog-library-directories:("." ".." "../or1200" "../jpeg" "../pkmc" "../dvga" "../uart" "../monitor" "../lab1" "../dafk_tb" "../eth" "../wb" "../leela")
// End:
