`include "include/timescale.v"

module or1200_vlx_su(/*AUTOARG*/
);

endmodule // or1200_vlx_su
// Local Variables:
// verilog-library-directories:("." ".." "../or1200" "../jpeg" "../pkmc" "../dvga" "../uart" "../monitor" "../lab1" "../dafk_tb" "../eth" "../wb" "../leela")
// End:
